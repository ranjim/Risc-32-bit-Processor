module programs (
    input clk,
    input en_read,
    input [31:0] pc,
    output reg [31:0] inst
);

parameter HALT = 0;
parameter NOP = 32'b00010000000000000000000000000000;

// define memory of 512 32-bit words
reg [31:0] mem [511:0];


initial begin
    mem[0] <= NOP;
    // store 10 numbers in registers 1-10 (R1-R10)
    // numbers are 11, 1, 67, 89, 69, 310, -12, 42, 0, 100
    mem[1] <= {3'b010, 3'b000, 16'b0000000000001011, 5'b00000, 5'b00001}; // R1 <- 11
    mem[2] <= {3'b010, 3'b000, 16'b0000000000000001, 5'b00000, 5'b00010}; // R2 <- 1
    mem[3] <= {3'b010, 3'b000, 16'b0000000001000011, 5'b00000, 5'b00011}; // R3 <- 67
    mem[4] <= {3'b010, 3'b000, 16'b0000000001011001, 5'b00000, 5'b00100}; // R4 <- 89
    mem[5] <= {3'b010, 3'b000, 16'b0000000001000101, 5'b00000, 5'b00101}; // R5 <- 69
    mem[6] <= {3'b010, 3'b000, 16'b0000000100110110, 5'b00000, 5'b00110}; // R6 <- 310
    mem[7] <= {3'b010, 3'b000, 16'b1111111111110100, 5'b00000, 5'b00111}; // R7 <- -12
    mem[8] <= {3'b010, 3'b000, 16'b0000000000101010, 5'b00000, 5'b01000}; // R8 <- 42
    mem[9] <= {3'b010, 3'b000, 16'b0000000000000000, 5'b00000, 5'b01001}; // R9 <- 0
    mem[10] <= {3'b010, 3'b000, 16'b0000000001100100, 5'b00000, 5'b01010}; // R10 <- 100
    mem[11] <= NOP;

    // now do bubble sort
    // do comparisons 45 times (10 choose 2)
    // each comparison is 3 instructions

    // first comparison
    mem[12] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    mem[13] <= {3'b101, 2'b10, 22'b0000000000000000010001, 5'b01111}; // if R15 > 0, jump to 17
    // swap R1 and R2 using R14 as temp
    mem[14] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[15] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[16] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[17] <= NOP;

    // second comparison
    mem[18] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    mem[19] <= {3'b101, 2'b10, 22'b0000000000000000010111, 5'b01111}; // if R15 > 0, jump to 23
    // swap R2 and R3 using R14 as temp
    mem[20] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[21] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[22] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[23] <= NOP;

    // third comparison
    mem[24] <= {3'b001, 3'b001, 11'b00000000000, 5'b00011, 5'b00100, 5'b01111}; // R4 - R3, store in R15
    mem[25] <= {3'b101, 2'b10, 22'b0000000000000000011101, 5'b01111}; // if R15 > 0, jump to 29
    // swap R3 and R4 using R14 as temp
    mem[26] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b01110}; // R14 <- R3
    mem[27] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b00011}; // R3 <- R4
    mem[28] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00100}; // R4 <- R14
    mem[29] <= NOP;

    // fourth comparison
    mem[30] <= {3'b001, 3'b001, 11'b00000000000, 5'b00100, 5'b00101, 5'b01111}; // R5 - R4, store in R15
    mem[31] <= {3'b101, 2'b10, 22'b0000000000000000100011, 5'b01111}; // if R15 > 0, jump to 35
    // swap R4 and R5 using R14 as temp
    mem[32] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b01110}; // R14 <- R4
    mem[33] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b00100}; // R4 <- R5
    mem[34] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00101}; // R5 <- R14
    mem[35] <= NOP;

    // fifth comparison
    mem[36] <= {3'b001, 3'b001, 11'b00000000000, 5'b00101, 5'b00110, 5'b01111}; // R6 - R5, store in R15
    mem[37] <= {3'b101, 2'b10, 22'b0000000000000000101001, 5'b01111}; // if R15 > 0, jump to 41
    // swap R5 and R6 using R14 as temp
    mem[38] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b01110}; // R14 <- R5
    mem[39] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b00101}; // R5 <- R6
    mem[40] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00110}; // R6 <- R14
    mem[41] <= NOP;

    // sixth comparison
    mem[42] <= {3'b001, 3'b001, 11'b00000000000, 5'b00110, 5'b00111, 5'b01111}; // R7 - R6, store in R15
    // if R15 > 0, jump to 47
    mem[43] <= {3'b101, 2'b10, 22'b0000000000000000101111, 5'b01111}; // if R15 > 0, jump to 47
    // swap R6 and R7 using R14 as temp
    mem[44] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b01110}; // R14 <- R6
    mem[45] <= {3'b111, 19'b0000000000000000000, 5'b00111, 5'b00110}; // R6 <- R7
    mem[46] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00111}; // R7 <- R14
    mem[47] <= NOP;

    // seventh comparison
    mem[48] <= {3'b001, 3'b001, 11'b00000000000, 5'b00111, 5'b01000, 5'b01111}; // R8 - R7, store in R15
    // if R15 > 0, jump to 53
    mem[49] <= {3'b101, 2'b10, 22'b0000000000000000110101, 5'b01111}; // if R15 > 0, jump to 53
    // swap R7 and R8 using R14 as temp
    mem[50] <= {3'b111, 19'b0000000000000000000, 5'b00111, 5'b01110}; // R14 <- R7
    mem[51] <= {3'b111, 19'b0000000000000000000, 5'b01000, 5'b00111}; // R7 <- R8
    mem[52] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b01000}; // R8 <- R14
    mem[53] <= NOP;

    // eighth comparison
    mem[54] <= {3'b001, 3'b001, 11'b00000000000, 5'b01000, 5'b01001, 5'b01111}; // R9 - R8, store in R15
    // if R15 > 0, jump to 59
    mem[55] <= {3'b101, 2'b10, 22'b0000000000000000111011, 5'b01111}; // if R15 > 0, jump to 59
    // swap R8 and R9 using R14 as temp
    mem[56] <= {3'b111, 19'b0000000000000000000, 5'b01000, 5'b01110}; // R14 <- R8
    mem[57] <= {3'b111, 19'b0000000000000000000, 5'b01001, 5'b01000}; // R8 <- R9
    mem[58] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b01001}; // R9 <- R14
    mem[59] <= NOP;

    // ninth comparison
    mem[60] <= {3'b001, 3'b001, 11'b00000000000, 5'b01001, 5'b01010, 5'b01111}; // R10 - R9, store in R15
    // if R15 > 0, jump to 65
    mem[61] <= {3'b101, 2'b10, 22'b0000000000000001000001, 5'b01111}; // if R15 > 0, jump to 65
    // swap R9 and R10 using R14 as temp
    mem[62] <= {3'b111, 19'b0000000000000000000, 5'b01001, 5'b01110}; // R14 <- R9
    mem[63] <= {3'b111, 19'b0000000000000000000, 5'b01010, 5'b01001}; // R9 <- R10
    mem[64] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b01010}; // R10 <- R14
    mem[65] <= NOP;

    // now largest number is in R10
    // repeat 9 times

    // tenth comparison
    mem[66] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 71
    mem[67] <= {3'b101, 2'b10, 22'b0000000000000001000111, 5'b01111}; // if R15 > 0, jump to 71
    // swap R1 and R2 using R14 as temp
    mem[68] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[69] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[70] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[71] <= NOP;

    // eleventh comparison
    mem[72] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    // if R15 > 0, jump to 77
    mem[73] <= {3'b101, 2'b10, 22'b0000000000000001001101, 5'b01111}; // if R15 > 0, jump to 77
    // swap R2 and R3 using R14 as temp
    mem[74] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[75] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[76] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[77] <= NOP;

    // twelfth comparison
    mem[78] <= {3'b001, 3'b001, 11'b00000000000, 5'b00011, 5'b00100, 5'b01111}; // R4 - R3, store in R15
    // if R15 > 0, jump to 83
    mem[79] <= {3'b101, 2'b10, 22'b0000000000000001010011, 5'b01111}; // if R15 > 0, jump to 83
    // swap R3 and R4 using R14 as temp
    mem[80] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b01110}; // R14 <- R3
    mem[81] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b00011}; // R3 <- R4
    mem[82] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00100}; // R4 <- R14
    mem[83] <= NOP;

    // thirteenth comparison
    mem[84] <= {3'b001, 3'b001, 11'b00000000000, 5'b00100, 5'b00101, 5'b01111}; // R5 - R4, store in R15
    // if R15 > 0, jump to 89
    mem[85] <= {3'b101, 2'b10, 22'b0000000000000001011001, 5'b01111}; // if R15 > 0, jump to 89
    // swap R4 and R5 using R14 as temp
    mem[86] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b01110}; // R14 <- R4
    mem[87] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b00100}; // R4 <- R5
    mem[88] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00101}; // R5 <- R14
    mem[89] <= NOP;

    // fourteenth comparison
    mem[90] <= {3'b001, 3'b001, 11'b00000000000, 5'b00101, 5'b00110, 5'b01111}; // R6 - R5, store in R15
    // if R15 > 0, jump to 95
    mem[91] <= {3'b101, 2'b10, 22'b0000000000000001011111, 5'b01111}; // if R15 > 0, jump to 95
    // swap R5 and R6 using R14 as temp
    mem[92] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b01110}; // R14 <- R5
    mem[93] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b00101}; // R5 <- R6
    mem[94] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00110}; // R6 <- R14
    mem[95] <= NOP;

    // fifteenth comparison
    mem[96] <= {3'b001, 3'b001, 11'b00000000000, 5'b00110, 5'b00111, 5'b01111}; // R7 - R6, store in R15
    // if R15 > 0, jump to 101
    mem[97] <= {3'b101, 2'b10, 22'b0000000000000001100101, 5'b01111}; // if R15 > 0, jump to 101
    // swap R6 and R7 using R14 as temp
    mem[98] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b01110}; // R14 <- R6
    mem[99] <= {3'b111, 19'b0000000000000000000, 5'b00111, 5'b00110}; // R6 <- R7
    mem[100] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00111}; // R7 <- R14
    mem[101] <= NOP;

    // sixteenth comparison
    mem[102] <= {3'b001, 3'b001, 11'b00000000000, 5'b00111, 5'b01000, 5'b01111}; // R8 - R7, store in R15
    // if R15 > 0, jump to 107
    mem[103] <= {3'b101, 2'b10, 22'b0000000000000001101011, 5'b01111}; // if R15 > 0, jump to 107
    // swap R7 and R8 using R14 as temp
    mem[104] <= {3'b111, 19'b0000000000000000000, 5'b00111, 5'b01110}; // R14 <- R7
    mem[105] <= {3'b111, 19'b0000000000000000000, 5'b01000, 5'b00111}; // R7 <- R8
    mem[106] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b01000}; // R8 <- R14
    mem[107] <= NOP;

    // seventeenth comparison
    mem[108] <= {3'b001, 3'b001, 11'b00000000000, 5'b01000, 5'b01001, 5'b01111}; // R9 - R8, store in R15
    // if R15 > 0, jump to 113
    mem[109] <= {3'b101, 2'b10, 22'b0000000000000001110001, 5'b01111}; // if R15 > 0, jump to 113
    // swap R8 and R9 using R14 as temp
    mem[110] <= {3'b111, 19'b0000000000000000000, 5'b01000, 5'b01110}; // R14 <- R8
    mem[111] <= {3'b111, 19'b0000000000000000000, 5'b01001, 5'b01000}; // R8 <- R9
    mem[112] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b01001}; // R9 <- R14
    mem[113] <= NOP;

    // now 2nd largest number is in R9
    // repeat 8 times

    // eighteenth comparison
    mem[114] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 119
    mem[115] <= {3'b101, 2'b10, 22'b0000000000000001110111, 5'b01111}; // if R15 > 0, jump to 119
    // swap R1 and R2 using R14 as temp
    mem[116] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[117] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[118] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[119] <= NOP;

    // nineteenth comparison
    mem[120] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    // if R15 > 0, jump to 125
    mem[121] <= {3'b101, 2'b10, 22'b0000000000000001111101, 5'b01111}; // if R15 > 0, jump to 125
    // swap R2 and R3 using R14 as temp
    mem[122] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[123] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[124] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[125] <= NOP;

    // twentieth comparison
    mem[126] <= {3'b001, 3'b001, 11'b00000000000, 5'b00011, 5'b00100, 5'b01111}; // R4 - R3, store in R15
    // if R15 > 0, jump to 131
    mem[127] <= {3'b101, 2'b10, 22'b0000000000000010000011, 5'b01111}; // if R15 > 0, jump to 131
    // swap R3 and R4 using R14 as temp
    mem[128] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b01110}; // R14 <- R3
    mem[129] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b00011}; // R3 <- R4
    mem[130] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00100}; // R4 <- R14
    mem[131] <= NOP;

    // twenty-first comparison
    mem[132] <= {3'b001, 3'b001, 11'b00000000000, 5'b00100, 5'b00101, 5'b01111}; // R5 - R4, store in R15
    // if R15 > 0, jump to 137
    mem[133] <= {3'b101, 2'b10, 22'b0000000000000010001001, 5'b01111}; // if R15 > 0, jump to 137
    // swap R4 and R5 using R14 as temp
    mem[134] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b01110}; // R14 <- R4
    mem[135] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b00100}; // R4 <- R5
    mem[136] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00101}; // R5 <- R14
    mem[137] <= NOP;

    // twenty-second comparison
    mem[138] <= {3'b001, 3'b001, 11'b00000000000, 5'b00101, 5'b00110, 5'b01111}; // R6 - R5, store in R15
    // if R15 > 0, jump to 143
    mem[139] <= {3'b101, 2'b10, 22'b0000000000000010001111, 5'b01111}; // if R15 > 0, jump to 143
    // swap R5 and R6 using R14 as temp
    mem[140] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b01110}; // R14 <- R5
    mem[141] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b00101}; // R5 <- R6
    mem[142] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00110}; // R6 <- R14
    mem[143] <= NOP;

    // twenty-third comparison
    mem[144] <= {3'b001, 3'b001, 11'b00000000000, 5'b00110, 5'b00111, 5'b01111}; // R7 - R6, store in R15
    // if R15 > 0, jump to 149
    mem[145] <= {3'b101, 2'b10, 22'b0000000000000010010101, 5'b01111}; // if R15 > 0, jump to 149
    // swap R6 and R7 using R14 as temp
    mem[146] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b01110}; // R14 <- R6
    mem[147] <= {3'b111, 19'b0000000000000000000, 5'b00111, 5'b00110}; // R6 <- R7
    mem[148] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00111}; // R7 <- R14
    mem[149] <= NOP;

    // twenty-fourth comparison
    mem[150] <= {3'b001, 3'b001, 11'b00000000000, 5'b00111, 5'b01000, 5'b01111}; // R8 - R7, store in R15
    // if R15 > 0, jump to 155
    mem[151] <= {3'b101, 2'b10, 22'b0000000000000010011011, 5'b01111}; // if R15 > 0, jump to 155
    // swap R7 and R8 using R14 as temp
    mem[152] <= {3'b111, 19'b0000000000000000000, 5'b00111, 5'b01110}; // R14 <- R7
    mem[153] <= {3'b111, 19'b0000000000000000000, 5'b01000, 5'b00111}; // R7 <- R8
    mem[154] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b01000}; // R8 <- R14
    mem[155] <= NOP;

    // now 3rd largest number is in R8
    // repeat 7 times

    // twenty-fifth comparison
    mem[156] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 161
    mem[157] <= {3'b101, 2'b10, 22'b0000000000000010100001, 5'b01111}; // if R15 > 0, jump to 161
    // swap R1 and R2 using R14 as temp
    mem[158] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[159] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[160] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[161] <= NOP;

    // twenty-sixth comparison
    mem[162] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    // if R15 > 0, jump to 167
    mem[163] <= {3'b101, 2'b10, 22'b0000000000000010100111, 5'b01111}; // if R15 > 0, jump to 167
    // swap R2 and R3 using R14 as temp
    mem[164] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[165] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[166] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[167] <= NOP;

    // twenty-seventh comparison
    mem[168] <= {3'b001, 3'b001, 11'b00000000000, 5'b00011, 5'b00100, 5'b01111}; // R4 - R3, store in R15
    // if R15 > 0, jump to 173
    mem[169] <= {3'b101, 2'b10, 22'b0000000000000010101101, 5'b01111}; // if R15 > 0, jump to 173
    // swap R3 and R4 using R14 as temp
    mem[170] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b01110}; // R14 <- R3
    mem[171] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b00011}; // R3 <- R4
    mem[172] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00100}; // R4 <- R14
    mem[173] <= NOP;

    // twenty-eighth comparison
    mem[174] <= {3'b001, 3'b001, 11'b00000000000, 5'b00100, 5'b00101, 5'b01111}; // R5 - R4, store in R15
    // if R15 > 0, jump to 179
    mem[175] <= {3'b101, 2'b10, 22'b0000000000000010110011, 5'b01111}; // if R15 > 0, jump to 179
    // swap R4 and R5 using R14 as temp
    mem[176] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b01110}; // R14 <- R4
    mem[177] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b00100}; // R4 <- R5
    mem[178] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00101}; // R5 <- R14
    mem[179] <= NOP;

    // twenty-ninth comparison
    mem[180] <= {3'b001, 3'b001, 11'b00000000000, 5'b00101, 5'b00110, 5'b01111}; // R6 - R5, store in R15
    // if R15 > 0, jump to 185
    mem[181] <= {3'b101, 2'b10, 22'b0000000000000010111001, 5'b01111}; // if R15 > 0, jump to 185
    // swap R5 and R6 using R14 as temp
    mem[182] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b01110}; // R14 <- R5
    mem[183] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b00101}; // R5 <- R6
    mem[184] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00110}; // R6 <- R14
    mem[185] <= NOP;

    // thirtieth comparison
    mem[186] <= {3'b001, 3'b001, 11'b00000000000, 5'b00110, 5'b00111, 5'b01111}; // R7 - R6, store in R15
    // if R15 > 0, jump to 191
    mem[187] <= {3'b101, 2'b10, 22'b0000000000000010111111, 5'b01111}; // if R15 > 0, jump to 191
    // swap R6 and R7 using R14 as temp
    mem[188] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b01110}; // R14 <- R6
    mem[189] <= {3'b111, 19'b0000000000000000000, 5'b00111, 5'b00110}; // R6 <- R7
    mem[190] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00111}; // R7 <- R14
    mem[191] <= NOP;

    // now 4th largest number is in R7
    // repeat 6 times

    // thirty-first comparison
    mem[192] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 197
    mem[193] <= {3'b101, 2'b10, 22'b0000000000000011000101, 5'b01111}; // if R15 > 0, jump to 197
    // swap R1 and R2 using R14 as temp
    mem[194] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[195] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[196] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[197] <= NOP;

    // thirty-second comparison
    mem[198] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    // if R15 > 0, jump to 203
    mem[199] <= {3'b101, 2'b10, 22'b0000000000000011001011, 5'b01111}; // if R15 > 0, jump to 203
    // swap R2 and R3 using R14 as temp
    mem[200] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[201] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[202] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[203] <= NOP;

    // thirty-third comparison
    mem[204] <= {3'b001, 3'b001, 11'b00000000000, 5'b00011, 5'b00100, 5'b01111}; // R4 - R3, store in R15
    // if R15 > 0, jump to 209
    mem[205] <= {3'b101, 2'b10, 22'b0000000000000011010001, 5'b01111}; // if R15 > 0, jump to 209
    // swap R3 and R4 using R14 as temp
    mem[206] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b01110}; // R14 <- R3
    mem[207] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b00011}; // R3 <- R4
    mem[208] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00100}; // R4 <- R14
    mem[209] <= NOP;

    // thirty-fourth comparison
    mem[210] <= {3'b001, 3'b001, 11'b00000000000, 5'b00100, 5'b00101, 5'b01111}; // R5 - R4, store in R15
    // if R15 > 0, jump to 215
    mem[211] <= {3'b101, 2'b10, 22'b0000000000000011010111, 5'b01111}; // if R15 > 0, jump to 215
    // swap R4 and R5 using R14 as temp
    mem[212] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b01110}; // R14 <- R4
    mem[213] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b00100}; // R4 <- R5
    mem[214] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00101}; // R5 <- R14
    mem[215] <= NOP;

    // thirty-fifth comparison
    mem[216] <= {3'b001, 3'b001, 11'b00000000000, 5'b00101, 5'b00110, 5'b01111}; // R6 - R5, store in R15
    // if R15 > 0, jump to 221
    mem[217] <= {3'b101, 2'b10, 22'b0000000000000011011101, 5'b01111}; // if R15 > 0, jump to 221
    // swap R5 and R6 using R14 as temp
    mem[218] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b01110}; // R14 <- R5
    mem[219] <= {3'b111, 19'b0000000000000000000, 5'b00110, 5'b00101}; // R5 <- R6
    mem[220] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00110}; // R6 <- R14
    mem[221] <= NOP;

    // now 5th largest number is in R6
    // repeat 5 times

    // thirty-sixth comparison
    mem[222] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 227
    mem[223] <= {3'b101, 2'b10, 22'b0000000000000011100011, 5'b01111}; // if R15 > 0, jump to 227
    // swap R1 and R2 using R14 as temp
    mem[224] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[225] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[226] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[227] <= NOP;

    // thirty-seventh comparison
    mem[228] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    // if R15 > 0, jump to 233
    mem[229] <= {3'b101, 2'b10, 22'b0000000000000011101001, 5'b01111}; // if R15 > 0, jump to 233
    // swap R2 and R3 using R14 as temp
    mem[230] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[231] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[232] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[233] <= NOP;

    // thirty-eighth comparison
    mem[234] <= {3'b001, 3'b001, 11'b00000000000, 5'b00011, 5'b00100, 5'b01111}; // R4 - R3, store in R15
    // if R15 > 0, jump to 239
    mem[235] <= {3'b101, 2'b10, 22'b0000000000000011101111, 5'b01111}; // if R15 > 0, jump to 239
    // swap R3 and R4 using R14 as temp
    mem[236] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b01110}; // R14 <- R3
    mem[237] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b00011}; // R3 <- R4
    mem[238] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00100}; // R4 <- R14
    mem[239] <= NOP;

    // thirty-ninth comparison
    mem[240] <= {3'b001, 3'b001, 11'b00000000000, 5'b00100, 5'b00101, 5'b01111}; // R5 - R4, store in R15
    // if R15 > 0, jump to 245
    mem[241] <= {3'b101, 2'b10, 22'b0000000000000011110101, 5'b01111}; // if R15 > 0, jump to 245
    // swap R4 and R5 using R14 as temp
    mem[242] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b01110}; // R14 <- R4
    mem[243] <= {3'b111, 19'b0000000000000000000, 5'b00101, 5'b00100}; // R4 <- R5
    mem[244] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00101}; // R5 <- R14
    mem[245] <= NOP;

    // now 6th largest number is in R5
    // repeat 4 times

    // fortieth comparison
    mem[246] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 251
    mem[247] <= {3'b101, 2'b10, 22'b0000000000000011111011, 5'b01111}; // if R15 > 0, jump to 251
    // swap R1 and R2 using R14 as temp
    mem[248] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[249] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[250] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[251] <= NOP;

    // forty-first comparison
    mem[252] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    // if R15 > 0, jump to 257
    mem[253] <= {3'b101, 2'b10, 22'b0000000000000100000001, 5'b01111}; // if R15 > 0, jump to 257
    // swap R2 and R3 using R14 as temp
    mem[254] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[255] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[256] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[257] <= NOP;

    // forty-second comparison
    mem[258] <= {3'b001, 3'b001, 11'b00000000000, 5'b00011, 5'b00100, 5'b01111}; // R4 - R3, store in R15
    // if R15 > 0, jump to 263
    mem[259] <= {3'b101, 2'b10, 22'b0000000000000100000111, 5'b01111}; // if R15 > 0, jump to 263
    // swap R3 and R4 using R14 as temp
    mem[260] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b01110}; // R14 <- R3
    mem[261] <= {3'b111, 19'b0000000000000000000, 5'b00100, 5'b00011}; // R3 <- R4
    mem[262] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00100}; // R4 <- R14
    mem[263] <= NOP;

    // now 7th largest number is in R4
    // repeat 3 times

    // forty-third comparison
    mem[264] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 269
    mem[265] <= {3'b101, 2'b10, 22'b0000000000000100001101, 5'b01111}; // if R15 > 0, jump to 269
    // swap R1 and R2 using R14 as temp
    mem[266] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[267] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[268] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[269] <= NOP;
    
    // forty-fourth comparison
    mem[270] <= {3'b001, 3'b001, 11'b00000000000, 5'b00010, 5'b00011, 5'b01111}; // R3 - R2, store in R15
    // if R15 > 0, jump to 275
    mem[271] <= {3'b101, 2'b10, 22'b0000000000000100010011, 5'b01111}; // if R15 > 0, jump to 275
    // swap R2 and R3 using R14 as temp
    mem[272] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b01110}; // R14 <- R2
    mem[273] <= {3'b111, 19'b0000000000000000000, 5'b00011, 5'b00010}; // R2 <- R3
    mem[274] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00011}; // R3 <- R14
    mem[275] <= NOP;

    // now 8th largest number is in R3
    // last comparison

    // forty-fifth comparison
    mem[276] <= {3'b001, 3'b001, 11'b00000000000, 5'b00001, 5'b00010, 5'b01111}; // R2 - R1, store in R15
    // if R15 > 0, jump to 281
    mem[277] <= {3'b101, 2'b10, 22'b0000000000000100011001, 5'b01111}; // if R15 > 0, jump to 281
    // swap R1 and R2 using R14 as temp
    mem[278] <= {3'b111, 19'b0000000000000000000, 5'b00001, 5'b01110}; // R14 <- R1
    mem[279] <= {3'b111, 19'b0000000000000000000, 5'b00010, 5'b00001}; // R1 <- R2
    mem[280] <= {3'b111, 19'b0000000000000000000, 5'b01110, 5'b00010}; // R2 <- R14
    mem[281] <= NOP;

    // now 9th largest number is in R2
    // smallest number is in R1

    mem[282] <= HALT;
end

always @(posedge clk) begin
    if (en_read) begin
        inst <= mem[pc];
    end
end

endmodule